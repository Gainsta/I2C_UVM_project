/*@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@|  File name   : i2c_pkg_inc.sv                                              @
@|  Project     : I2C_Test :: I2C                                            @
@|  Created     : Nikolay Dvoynishnikov                                     @
@|  Description : Include packages for I2C testbench                        @
@|  Data        :  - .12.2020                                                @
@|  Notes                                                                     @
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@*/

`ifndef I2C_PACKAGE_INC__
`define I2C_PACKAGE_INC__

//------------------------------------------------------
// UVM package
`include "uvm_pkg.sv"

`endif // I2C_PACKAGE_INC__